module CheckAlg(
	
	input logic qb,
	output logic flag

);

	always_comb
	begin
		if (qb == 1) begin
			flag = 1;
		end
	end
endmodule
