module logic_Module
(
	input logic up_state,        
	input logic down_state,
	input logic left_state,
	input logic right_state,
	output logic lose_output,
	output logic win_output,
	
	output logic [15:0][3:0] cell_matrix
	
	//input logic clk (????)   
	
);




endmodule