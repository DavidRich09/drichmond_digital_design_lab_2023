//module countdown_nbits_tb;
//
//
//parameter CLK = 10; 
//
//reg clk;
//reg rst;
//wire [N-1:0] countdownOut;
//
//
//countdown_timer dut (
//  .clk(clk),
//  .rst(rst),
//  .countdownOut(countdownOut)
//);
//
//
//initial begin
//
//// test 2 bits
//
//
//
//
//
//
//
//
//end
//
//endmodule