module ALU 	

(
);



endmodule