module Control_Unit_Decoder 	

(
	input logic [1:0] op,        
	input logic [5:0] funct,
	input logic [3:0] rd,
	output logic pcs,
	output logic reg_w,
	output logic mem_w,
	output logic mem_to_reg,
	output logic alu_src,
	output logic [1:0] flag_w,
	output logic [1:0] imm_src,
	output logic [1:0] reg_src,
	output logic [1:0] alu_control

);



endmodule