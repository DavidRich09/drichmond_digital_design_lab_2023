module control_unit_tb;

   // Señales del test bench


   // Instancia del módulo bajo prueba


   initial begin
	
   end


endmodule