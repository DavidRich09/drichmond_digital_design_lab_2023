module Processor_Image 	

(
   

);



endmodule