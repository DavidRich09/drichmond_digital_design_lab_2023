module VGA_Main_Module
(

	input logic [15:0][3:0] cell_matrix
	
	//output logic ????? @Sergio ahí ve que hace
	 
);




endmodule