module maquina_Estados

(
	input logic up,        
	input logic down,
	input logic left,
	input logic right,
	input logic logic_lose_input,
	input logic logic_win_input,
	
	output logic up_state,        
	output logic down_state,
	output logic left_state,
	output logic right_state
	//output logic lose_state,
	//output logic win_state
	
	//input logic clk (????)   
	
);




endmodule